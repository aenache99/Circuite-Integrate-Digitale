module tb();
reg instruction_tb;
reg data0_tb;
reg data1_tb;
wire overflow_flag_tb;
wire zero_flag;
wire out0_tb;
wire out1_tb;
wire out2_tb;
wire out3_tb;
// instantiere DUT:
top DUT(.instruction(instruction_tb),
			.data0(data0_tb),
			.data1(data1_tb),
			.overflow_flag(overflow_flag_tb),
			.zero_flag(zero_flag_tb),
			.out0(out0_tb),
			.out1(out1_tb),
			.out2(out2_tb),
			.out3(out3_tb));
//Dam valori:
initial
begin
	instruction_tb = 0;
	data0_tb = 0;
	data1_tb = 0;
	#10 instruction_tb = 16'hffff;
	#20 data0_tb = 255;
		data1_tb = 255;
	#30 instruction_tb = 16'b00_00_10_00000000;
		data0_tb = 1;
		data1_tb = 1;
	#35 data0_tb = 2;
	#40 data1_tb = 3;
end
// Oprire simulare:
initial 
begin
	#1000 $stop;
end
endmodule

// n-am mai avut timp sa ma uit in modelsim, rip me :(
