module ParityChecker(input wire [3:0]in,
							output wire out
							);

assign out = in[0];
endmodule 