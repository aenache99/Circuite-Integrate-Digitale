module sumator(input [2:0] in0,
					input [2:0] in1,
					output [3:0] out
);
assign out=in0+in1;
endmodule 