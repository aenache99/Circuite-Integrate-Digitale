module not_gate (
				input wire in0,
				output wire out0
				);
				
assign out0 = !in0;
endmodule //not_gate