module mux44bit(input wire [3:0]in0,
				  input wire [3:0]in1,
				  input wire [3:0]in2,
				  input wire [3:0]in3,
				  input wire [1:0]sel,
				  output wire [3:0]out
				  );
assign out = sel[1] ? (sel[0] ? in3 : in2) : (sel[0] ? in1 : in0);
endmodule 